module layer0 (input [127:0] M0, output [255:0] M1);

wire [7:0] layer0_N0_wire = {M0[93], M0[92], M0[89], M0[88], M0[35], M0[34], M0[7], M0[6]};
layer0_N0 layer0_N0_inst (.M0(layer0_N0_wire), .M1(M1[1:0]));

wire [7:0] layer0_N1_wire = {M0[101], M0[100], M0[51], M0[50], M0[47], M0[46], M0[17], M0[16]};
layer0_N1 layer0_N1_inst (.M0(layer0_N1_wire), .M1(M1[3:2]));

wire [7:0] layer0_N2_wire = {M0[125], M0[124], M0[99], M0[98], M0[71], M0[70], M0[41], M0[40]};
layer0_N2 layer0_N2_inst (.M0(layer0_N2_wire), .M1(M1[5:4]));

wire [7:0] layer0_N3_wire = {M0[117], M0[116], M0[77], M0[76], M0[55], M0[54], M0[9], M0[8]};
layer0_N3 layer0_N3_inst (.M0(layer0_N3_wire), .M1(M1[7:6]));

wire [7:0] layer0_N4_wire = {M0[115], M0[114], M0[81], M0[80], M0[45], M0[44], M0[19], M0[18]};
layer0_N4 layer0_N4_inst (.M0(layer0_N4_wire), .M1(M1[9:8]));

wire [7:0] layer0_N5_wire = {M0[67], M0[66], M0[51], M0[50], M0[49], M0[48], M0[7], M0[6]};
layer0_N5 layer0_N5_inst (.M0(layer0_N5_wire), .M1(M1[11:10]));

wire [7:0] layer0_N6_wire = {M0[75], M0[74], M0[57], M0[56], M0[37], M0[36], M0[35], M0[34]};
layer0_N6 layer0_N6_inst (.M0(layer0_N6_wire), .M1(M1[13:12]));

wire [7:0] layer0_N7_wire = {M0[101], M0[100], M0[65], M0[64], M0[39], M0[38], M0[15], M0[14]};
layer0_N7 layer0_N7_inst (.M0(layer0_N7_wire), .M1(M1[15:14]));

wire [7:0] layer0_N8_wire = {M0[123], M0[122], M0[119], M0[118], M0[93], M0[92], M0[37], M0[36]};
layer0_N8 layer0_N8_inst (.M0(layer0_N8_wire), .M1(M1[17:16]));

wire [7:0] layer0_N9_wire = {M0[103], M0[102], M0[81], M0[80], M0[59], M0[58], M0[37], M0[36]};
layer0_N9 layer0_N9_inst (.M0(layer0_N9_wire), .M1(M1[19:18]));

wire [7:0] layer0_N10_wire = {M0[117], M0[116], M0[113], M0[112], M0[45], M0[44], M0[35], M0[34]};
layer0_N10 layer0_N10_inst (.M0(layer0_N10_wire), .M1(M1[21:20]));

wire [7:0] layer0_N11_wire = {M0[95], M0[94], M0[75], M0[74], M0[69], M0[68], M0[65], M0[64]};
layer0_N11 layer0_N11_inst (.M0(layer0_N11_wire), .M1(M1[23:22]));

wire [7:0] layer0_N12_wire = {M0[103], M0[102], M0[91], M0[90], M0[75], M0[74], M0[13], M0[12]};
layer0_N12 layer0_N12_inst (.M0(layer0_N12_wire), .M1(M1[25:24]));

wire [7:0] layer0_N13_wire = {M0[125], M0[124], M0[55], M0[54], M0[45], M0[44], M0[5], M0[4]};
layer0_N13 layer0_N13_inst (.M0(layer0_N13_wire), .M1(M1[27:26]));

wire [7:0] layer0_N14_wire = {M0[95], M0[94], M0[45], M0[44], M0[39], M0[38], M0[35], M0[34]};
layer0_N14 layer0_N14_inst (.M0(layer0_N14_wire), .M1(M1[29:28]));

wire [7:0] layer0_N15_wire = {M0[109], M0[108], M0[77], M0[76], M0[53], M0[52], M0[45], M0[44]};
layer0_N15 layer0_N15_inst (.M0(layer0_N15_wire), .M1(M1[31:30]));

wire [7:0] layer0_N16_wire = {M0[85], M0[84], M0[45], M0[44], M0[39], M0[38], M0[29], M0[28]};
layer0_N16 layer0_N16_inst (.M0(layer0_N16_wire), .M1(M1[33:32]));

wire [7:0] layer0_N17_wire = {M0[91], M0[90], M0[55], M0[54], M0[41], M0[40], M0[25], M0[24]};
layer0_N17 layer0_N17_inst (.M0(layer0_N17_wire), .M1(M1[35:34]));

wire [7:0] layer0_N18_wire = {M0[111], M0[110], M0[79], M0[78], M0[41], M0[40], M0[7], M0[6]};
layer0_N18 layer0_N18_inst (.M0(layer0_N18_wire), .M1(M1[37:36]));

wire [7:0] layer0_N19_wire = {M0[99], M0[98], M0[65], M0[64], M0[35], M0[34], M0[3], M0[2]};
layer0_N19 layer0_N19_inst (.M0(layer0_N19_wire), .M1(M1[39:38]));

wire [7:0] layer0_N20_wire = {M0[123], M0[122], M0[109], M0[108], M0[75], M0[74], M0[31], M0[30]};
layer0_N20 layer0_N20_inst (.M0(layer0_N20_wire), .M1(M1[41:40]));

wire [7:0] layer0_N21_wire = {M0[109], M0[108], M0[41], M0[40], M0[35], M0[34], M0[5], M0[4]};
layer0_N21 layer0_N21_inst (.M0(layer0_N21_wire), .M1(M1[43:42]));

wire [7:0] layer0_N22_wire = {M0[99], M0[98], M0[57], M0[56], M0[53], M0[52], M0[47], M0[46]};
layer0_N22 layer0_N22_inst (.M0(layer0_N22_wire), .M1(M1[45:44]));

wire [7:0] layer0_N23_wire = {M0[99], M0[98], M0[69], M0[68], M0[25], M0[24], M0[1], M0[0]};
layer0_N23 layer0_N23_inst (.M0(layer0_N23_wire), .M1(M1[47:46]));

wire [7:0] layer0_N24_wire = {M0[115], M0[114], M0[113], M0[112], M0[13], M0[12], M0[3], M0[2]};
layer0_N24 layer0_N24_inst (.M0(layer0_N24_wire), .M1(M1[49:48]));

wire [7:0] layer0_N25_wire = {M0[63], M0[62], M0[55], M0[54], M0[47], M0[46], M0[29], M0[28]};
layer0_N25 layer0_N25_inst (.M0(layer0_N25_wire), .M1(M1[51:50]));

wire [7:0] layer0_N26_wire = {M0[49], M0[48], M0[43], M0[42], M0[27], M0[26], M0[17], M0[16]};
layer0_N26 layer0_N26_inst (.M0(layer0_N26_wire), .M1(M1[53:52]));

wire [7:0] layer0_N27_wire = {M0[121], M0[120], M0[109], M0[108], M0[95], M0[94], M0[77], M0[76]};
layer0_N27 layer0_N27_inst (.M0(layer0_N27_wire), .M1(M1[55:54]));

wire [7:0] layer0_N28_wire = {M0[105], M0[104], M0[95], M0[94], M0[85], M0[84], M0[1], M0[0]};
layer0_N28 layer0_N28_inst (.M0(layer0_N28_wire), .M1(M1[57:56]));

wire [7:0] layer0_N29_wire = {M0[55], M0[54], M0[45], M0[44], M0[31], M0[30], M0[15], M0[14]};
layer0_N29 layer0_N29_inst (.M0(layer0_N29_wire), .M1(M1[59:58]));

wire [7:0] layer0_N30_wire = {M0[109], M0[108], M0[107], M0[106], M0[85], M0[84], M0[67], M0[66]};
layer0_N30 layer0_N30_inst (.M0(layer0_N30_wire), .M1(M1[61:60]));

wire [7:0] layer0_N31_wire = {M0[61], M0[60], M0[31], M0[30], M0[21], M0[20], M0[5], M0[4]};
layer0_N31 layer0_N31_inst (.M0(layer0_N31_wire), .M1(M1[63:62]));

wire [7:0] layer0_N32_wire = {M0[119], M0[118], M0[65], M0[64], M0[15], M0[14], M0[11], M0[10]};
layer0_N32 layer0_N32_inst (.M0(layer0_N32_wire), .M1(M1[65:64]));

wire [7:0] layer0_N33_wire = {M0[113], M0[112], M0[47], M0[46], M0[45], M0[44], M0[5], M0[4]};
layer0_N33 layer0_N33_inst (.M0(layer0_N33_wire), .M1(M1[67:66]));

wire [7:0] layer0_N34_wire = {M0[127], M0[126], M0[113], M0[112], M0[95], M0[94], M0[9], M0[8]};
layer0_N34 layer0_N34_inst (.M0(layer0_N34_wire), .M1(M1[69:68]));

wire [7:0] layer0_N35_wire = {M0[85], M0[84], M0[71], M0[70], M0[57], M0[56], M0[49], M0[48]};
layer0_N35 layer0_N35_inst (.M0(layer0_N35_wire), .M1(M1[71:70]));

wire [7:0] layer0_N36_wire = {M0[115], M0[114], M0[93], M0[92], M0[47], M0[46], M0[15], M0[14]};
layer0_N36 layer0_N36_inst (.M0(layer0_N36_wire), .M1(M1[73:72]));

wire [7:0] layer0_N37_wire = {M0[87], M0[86], M0[71], M0[70], M0[67], M0[66], M0[25], M0[24]};
layer0_N37 layer0_N37_inst (.M0(layer0_N37_wire), .M1(M1[75:74]));

wire [7:0] layer0_N38_wire = {M0[125], M0[124], M0[121], M0[120], M0[105], M0[104], M0[81], M0[80]};
layer0_N38 layer0_N38_inst (.M0(layer0_N38_wire), .M1(M1[77:76]));

wire [7:0] layer0_N39_wire = {M0[117], M0[116], M0[93], M0[92], M0[39], M0[38], M0[37], M0[36]};
layer0_N39 layer0_N39_inst (.M0(layer0_N39_wire), .M1(M1[79:78]));

wire [7:0] layer0_N40_wire = {M0[127], M0[126], M0[113], M0[112], M0[105], M0[104], M0[53], M0[52]};
layer0_N40 layer0_N40_inst (.M0(layer0_N40_wire), .M1(M1[81:80]));

wire [7:0] layer0_N41_wire = {M0[125], M0[124], M0[113], M0[112], M0[85], M0[84], M0[79], M0[78]};
layer0_N41 layer0_N41_inst (.M0(layer0_N41_wire), .M1(M1[83:82]));

wire [7:0] layer0_N42_wire = {M0[117], M0[116], M0[75], M0[74], M0[69], M0[68], M0[47], M0[46]};
layer0_N42 layer0_N42_inst (.M0(layer0_N42_wire), .M1(M1[85:84]));

wire [7:0] layer0_N43_wire = {M0[109], M0[108], M0[75], M0[74], M0[65], M0[64], M0[9], M0[8]};
layer0_N43 layer0_N43_inst (.M0(layer0_N43_wire), .M1(M1[87:86]));

wire [7:0] layer0_N44_wire = {M0[119], M0[118], M0[79], M0[78], M0[13], M0[12], M0[9], M0[8]};
layer0_N44 layer0_N44_inst (.M0(layer0_N44_wire), .M1(M1[89:88]));

wire [7:0] layer0_N45_wire = {M0[119], M0[118], M0[107], M0[106], M0[59], M0[58], M0[1], M0[0]};
layer0_N45 layer0_N45_inst (.M0(layer0_N45_wire), .M1(M1[91:90]));

wire [7:0] layer0_N46_wire = {M0[113], M0[112], M0[47], M0[46], M0[43], M0[42], M0[17], M0[16]};
layer0_N46 layer0_N46_inst (.M0(layer0_N46_wire), .M1(M1[93:92]));

wire [7:0] layer0_N47_wire = {M0[113], M0[112], M0[99], M0[98], M0[23], M0[22], M0[17], M0[16]};
layer0_N47 layer0_N47_inst (.M0(layer0_N47_wire), .M1(M1[95:94]));

wire [7:0] layer0_N48_wire = {M0[89], M0[88], M0[59], M0[58], M0[41], M0[40], M0[17], M0[16]};
layer0_N48 layer0_N48_inst (.M0(layer0_N48_wire), .M1(M1[97:96]));

wire [7:0] layer0_N49_wire = {M0[107], M0[106], M0[53], M0[52], M0[49], M0[48], M0[45], M0[44]};
layer0_N49 layer0_N49_inst (.M0(layer0_N49_wire), .M1(M1[99:98]));

wire [7:0] layer0_N50_wire = {M0[81], M0[80], M0[63], M0[62], M0[21], M0[20], M0[5], M0[4]};
layer0_N50 layer0_N50_inst (.M0(layer0_N50_wire), .M1(M1[101:100]));

wire [7:0] layer0_N51_wire = {M0[103], M0[102], M0[99], M0[98], M0[31], M0[30], M0[17], M0[16]};
layer0_N51 layer0_N51_inst (.M0(layer0_N51_wire), .M1(M1[103:102]));

wire [7:0] layer0_N52_wire = {M0[89], M0[88], M0[87], M0[86], M0[69], M0[68], M0[11], M0[10]};
layer0_N52 layer0_N52_inst (.M0(layer0_N52_wire), .M1(M1[105:104]));

wire [7:0] layer0_N53_wire = {M0[125], M0[124], M0[101], M0[100], M0[17], M0[16], M0[5], M0[4]};
layer0_N53 layer0_N53_inst (.M0(layer0_N53_wire), .M1(M1[107:106]));

wire [7:0] layer0_N54_wire = {M0[111], M0[110], M0[93], M0[92], M0[73], M0[72], M0[15], M0[14]};
layer0_N54 layer0_N54_inst (.M0(layer0_N54_wire), .M1(M1[109:108]));

wire [7:0] layer0_N55_wire = {M0[97], M0[96], M0[75], M0[74], M0[47], M0[46], M0[31], M0[30]};
layer0_N55 layer0_N55_inst (.M0(layer0_N55_wire), .M1(M1[111:110]));

wire [7:0] layer0_N56_wire = {M0[33], M0[32], M0[21], M0[20], M0[19], M0[18], M0[11], M0[10]};
layer0_N56 layer0_N56_inst (.M0(layer0_N56_wire), .M1(M1[113:112]));

wire [7:0] layer0_N57_wire = {M0[125], M0[124], M0[73], M0[72], M0[27], M0[26], M0[21], M0[20]};
layer0_N57 layer0_N57_inst (.M0(layer0_N57_wire), .M1(M1[115:114]));

wire [7:0] layer0_N58_wire = {M0[115], M0[114], M0[103], M0[102], M0[95], M0[94], M0[3], M0[2]};
layer0_N58 layer0_N58_inst (.M0(layer0_N58_wire), .M1(M1[117:116]));

wire [7:0] layer0_N59_wire = {M0[55], M0[54], M0[41], M0[40], M0[35], M0[34], M0[17], M0[16]};
layer0_N59 layer0_N59_inst (.M0(layer0_N59_wire), .M1(M1[119:118]));

wire [7:0] layer0_N60_wire = {M0[89], M0[88], M0[53], M0[52], M0[5], M0[4], M0[3], M0[2]};
layer0_N60 layer0_N60_inst (.M0(layer0_N60_wire), .M1(M1[121:120]));

wire [7:0] layer0_N61_wire = {M0[81], M0[80], M0[77], M0[76], M0[75], M0[74], M0[19], M0[18]};
layer0_N61 layer0_N61_inst (.M0(layer0_N61_wire), .M1(M1[123:122]));

wire [7:0] layer0_N62_wire = {M0[127], M0[126], M0[93], M0[92], M0[81], M0[80], M0[37], M0[36]};
layer0_N62 layer0_N62_inst (.M0(layer0_N62_wire), .M1(M1[125:124]));

wire [7:0] layer0_N63_wire = {M0[117], M0[116], M0[115], M0[114], M0[107], M0[106], M0[85], M0[84]};
layer0_N63 layer0_N63_inst (.M0(layer0_N63_wire), .M1(M1[127:126]));

wire [7:0] layer0_N64_wire = {M0[121], M0[120], M0[119], M0[118], M0[99], M0[98], M0[69], M0[68]};
layer0_N64 layer0_N64_inst (.M0(layer0_N64_wire), .M1(M1[129:128]));

wire [7:0] layer0_N65_wire = {M0[61], M0[60], M0[43], M0[42], M0[35], M0[34], M0[21], M0[20]};
layer0_N65 layer0_N65_inst (.M0(layer0_N65_wire), .M1(M1[131:130]));

wire [7:0] layer0_N66_wire = {M0[117], M0[116], M0[111], M0[110], M0[97], M0[96], M0[61], M0[60]};
layer0_N66 layer0_N66_inst (.M0(layer0_N66_wire), .M1(M1[133:132]));

wire [7:0] layer0_N67_wire = {M0[121], M0[120], M0[117], M0[116], M0[25], M0[24], M0[5], M0[4]};
layer0_N67 layer0_N67_inst (.M0(layer0_N67_wire), .M1(M1[135:134]));

wire [7:0] layer0_N68_wire = {M0[67], M0[66], M0[37], M0[36], M0[21], M0[20], M0[7], M0[6]};
layer0_N68 layer0_N68_inst (.M0(layer0_N68_wire), .M1(M1[137:136]));

wire [7:0] layer0_N69_wire = {M0[97], M0[96], M0[71], M0[70], M0[53], M0[52], M0[39], M0[38]};
layer0_N69 layer0_N69_inst (.M0(layer0_N69_wire), .M1(M1[139:138]));

wire [7:0] layer0_N70_wire = {M0[105], M0[104], M0[71], M0[70], M0[69], M0[68], M0[5], M0[4]};
layer0_N70 layer0_N70_inst (.M0(layer0_N70_wire), .M1(M1[141:140]));

wire [7:0] layer0_N71_wire = {M0[93], M0[92], M0[77], M0[76], M0[75], M0[74], M0[69], M0[68]};
layer0_N71 layer0_N71_inst (.M0(layer0_N71_wire), .M1(M1[143:142]));

wire [7:0] layer0_N72_wire = {M0[101], M0[100], M0[95], M0[94], M0[89], M0[88], M0[81], M0[80]};
layer0_N72 layer0_N72_inst (.M0(layer0_N72_wire), .M1(M1[145:144]));

wire [7:0] layer0_N73_wire = {M0[101], M0[100], M0[79], M0[78], M0[41], M0[40], M0[21], M0[20]};
layer0_N73 layer0_N73_inst (.M0(layer0_N73_wire), .M1(M1[147:146]));

wire [7:0] layer0_N74_wire = {M0[53], M0[52], M0[39], M0[38], M0[37], M0[36], M0[33], M0[32]};
layer0_N74 layer0_N74_inst (.M0(layer0_N74_wire), .M1(M1[149:148]));

wire [7:0] layer0_N75_wire = {M0[25], M0[24], M0[19], M0[18], M0[15], M0[14], M0[11], M0[10]};
layer0_N75 layer0_N75_inst (.M0(layer0_N75_wire), .M1(M1[151:150]));

wire [7:0] layer0_N76_wire = {M0[121], M0[120], M0[107], M0[106], M0[25], M0[24], M0[3], M0[2]};
layer0_N76 layer0_N76_inst (.M0(layer0_N76_wire), .M1(M1[153:152]));

wire [7:0] layer0_N77_wire = {M0[123], M0[122], M0[101], M0[100], M0[69], M0[68], M0[19], M0[18]};
layer0_N77 layer0_N77_inst (.M0(layer0_N77_wire), .M1(M1[155:154]));

wire [7:0] layer0_N78_wire = {M0[69], M0[68], M0[57], M0[56], M0[19], M0[18], M0[5], M0[4]};
layer0_N78 layer0_N78_inst (.M0(layer0_N78_wire), .M1(M1[157:156]));

wire [7:0] layer0_N79_wire = {M0[95], M0[94], M0[57], M0[56], M0[17], M0[16], M0[1], M0[0]};
layer0_N79 layer0_N79_inst (.M0(layer0_N79_wire), .M1(M1[159:158]));

wire [7:0] layer0_N80_wire = {M0[99], M0[98], M0[35], M0[34], M0[25], M0[24], M0[9], M0[8]};
layer0_N80 layer0_N80_inst (.M0(layer0_N80_wire), .M1(M1[161:160]));

wire [7:0] layer0_N81_wire = {M0[127], M0[126], M0[125], M0[124], M0[89], M0[88], M0[35], M0[34]};
layer0_N81 layer0_N81_inst (.M0(layer0_N81_wire), .M1(M1[163:162]));

wire [7:0] layer0_N82_wire = {M0[99], M0[98], M0[93], M0[92], M0[85], M0[84], M0[17], M0[16]};
layer0_N82 layer0_N82_inst (.M0(layer0_N82_wire), .M1(M1[165:164]));

wire [7:0] layer0_N83_wire = {M0[125], M0[124], M0[117], M0[116], M0[73], M0[72], M0[9], M0[8]};
layer0_N83 layer0_N83_inst (.M0(layer0_N83_wire), .M1(M1[167:166]));

wire [7:0] layer0_N84_wire = {M0[113], M0[112], M0[81], M0[80], M0[77], M0[76], M0[53], M0[52]};
layer0_N84 layer0_N84_inst (.M0(layer0_N84_wire), .M1(M1[169:168]));

wire [7:0] layer0_N85_wire = {M0[119], M0[118], M0[105], M0[104], M0[97], M0[96], M0[93], M0[92]};
layer0_N85 layer0_N85_inst (.M0(layer0_N85_wire), .M1(M1[171:170]));

wire [7:0] layer0_N86_wire = {M0[71], M0[70], M0[23], M0[22], M0[19], M0[18], M0[5], M0[4]};
layer0_N86 layer0_N86_inst (.M0(layer0_N86_wire), .M1(M1[173:172]));

wire [7:0] layer0_N87_wire = {M0[93], M0[92], M0[91], M0[90], M0[89], M0[88], M0[63], M0[62]};
layer0_N87 layer0_N87_inst (.M0(layer0_N87_wire), .M1(M1[175:174]));

wire [7:0] layer0_N88_wire = {M0[91], M0[90], M0[87], M0[86], M0[69], M0[68], M0[5], M0[4]};
layer0_N88 layer0_N88_inst (.M0(layer0_N88_wire), .M1(M1[177:176]));

wire [7:0] layer0_N89_wire = {M0[107], M0[106], M0[89], M0[88], M0[57], M0[56], M0[37], M0[36]};
layer0_N89 layer0_N89_inst (.M0(layer0_N89_wire), .M1(M1[179:178]));

wire [7:0] layer0_N90_wire = {M0[115], M0[114], M0[83], M0[82], M0[37], M0[36], M0[1], M0[0]};
layer0_N90 layer0_N90_inst (.M0(layer0_N90_wire), .M1(M1[181:180]));

wire [7:0] layer0_N91_wire = {M0[105], M0[104], M0[91], M0[90], M0[49], M0[48], M0[11], M0[10]};
layer0_N91 layer0_N91_inst (.M0(layer0_N91_wire), .M1(M1[183:182]));

wire [7:0] layer0_N92_wire = {M0[121], M0[120], M0[89], M0[88], M0[43], M0[42], M0[17], M0[16]};
layer0_N92 layer0_N92_inst (.M0(layer0_N92_wire), .M1(M1[185:184]));

wire [7:0] layer0_N93_wire = {M0[113], M0[112], M0[79], M0[78], M0[53], M0[52], M0[31], M0[30]};
layer0_N93 layer0_N93_inst (.M0(layer0_N93_wire), .M1(M1[187:186]));

wire [7:0] layer0_N94_wire = {M0[87], M0[86], M0[61], M0[60], M0[43], M0[42], M0[5], M0[4]};
layer0_N94 layer0_N94_inst (.M0(layer0_N94_wire), .M1(M1[189:188]));

wire [7:0] layer0_N95_wire = {M0[105], M0[104], M0[97], M0[96], M0[93], M0[92], M0[59], M0[58]};
layer0_N95 layer0_N95_inst (.M0(layer0_N95_wire), .M1(M1[191:190]));

wire [7:0] layer0_N96_wire = {M0[85], M0[84], M0[59], M0[58], M0[21], M0[20], M0[11], M0[10]};
layer0_N96 layer0_N96_inst (.M0(layer0_N96_wire), .M1(M1[193:192]));

wire [7:0] layer0_N97_wire = {M0[103], M0[102], M0[57], M0[56], M0[49], M0[48], M0[9], M0[8]};
layer0_N97 layer0_N97_inst (.M0(layer0_N97_wire), .M1(M1[195:194]));

wire [7:0] layer0_N98_wire = {M0[101], M0[100], M0[93], M0[92], M0[79], M0[78], M0[23], M0[22]};
layer0_N98 layer0_N98_inst (.M0(layer0_N98_wire), .M1(M1[197:196]));

wire [7:0] layer0_N99_wire = {M0[75], M0[74], M0[63], M0[62], M0[19], M0[18], M0[7], M0[6]};
layer0_N99 layer0_N99_inst (.M0(layer0_N99_wire), .M1(M1[199:198]));

wire [7:0] layer0_N100_wire = {M0[81], M0[80], M0[67], M0[66], M0[41], M0[40], M0[25], M0[24]};
layer0_N100 layer0_N100_inst (.M0(layer0_N100_wire), .M1(M1[201:200]));

wire [7:0] layer0_N101_wire = {M0[99], M0[98], M0[79], M0[78], M0[37], M0[36], M0[29], M0[28]};
layer0_N101 layer0_N101_inst (.M0(layer0_N101_wire), .M1(M1[203:202]));

wire [7:0] layer0_N102_wire = {M0[121], M0[120], M0[115], M0[114], M0[109], M0[108], M0[15], M0[14]};
layer0_N102 layer0_N102_inst (.M0(layer0_N102_wire), .M1(M1[205:204]));

wire [7:0] layer0_N103_wire = {M0[117], M0[116], M0[83], M0[82], M0[75], M0[74], M0[67], M0[66]};
layer0_N103 layer0_N103_inst (.M0(layer0_N103_wire), .M1(M1[207:206]));

wire [7:0] layer0_N104_wire = {M0[127], M0[126], M0[67], M0[66], M0[35], M0[34], M0[3], M0[2]};
layer0_N104 layer0_N104_inst (.M0(layer0_N104_wire), .M1(M1[209:208]));

wire [7:0] layer0_N105_wire = {M0[125], M0[124], M0[47], M0[46], M0[23], M0[22], M0[17], M0[16]};
layer0_N105 layer0_N105_inst (.M0(layer0_N105_wire), .M1(M1[211:210]));

wire [7:0] layer0_N106_wire = {M0[79], M0[78], M0[19], M0[18], M0[9], M0[8], M0[3], M0[2]};
layer0_N106 layer0_N106_inst (.M0(layer0_N106_wire), .M1(M1[213:212]));

wire [7:0] layer0_N107_wire = {M0[115], M0[114], M0[101], M0[100], M0[75], M0[74], M0[53], M0[52]};
layer0_N107 layer0_N107_inst (.M0(layer0_N107_wire), .M1(M1[215:214]));

wire [7:0] layer0_N108_wire = {M0[119], M0[118], M0[81], M0[80], M0[75], M0[74], M0[69], M0[68]};
layer0_N108 layer0_N108_inst (.M0(layer0_N108_wire), .M1(M1[217:216]));

wire [7:0] layer0_N109_wire = {M0[117], M0[116], M0[91], M0[90], M0[45], M0[44], M0[35], M0[34]};
layer0_N109 layer0_N109_inst (.M0(layer0_N109_wire), .M1(M1[219:218]));

wire [7:0] layer0_N110_wire = {M0[121], M0[120], M0[115], M0[114], M0[85], M0[84], M0[1], M0[0]};
layer0_N110 layer0_N110_inst (.M0(layer0_N110_wire), .M1(M1[221:220]));

wire [7:0] layer0_N111_wire = {M0[115], M0[114], M0[73], M0[72], M0[71], M0[70], M0[7], M0[6]};
layer0_N111 layer0_N111_inst (.M0(layer0_N111_wire), .M1(M1[223:222]));

wire [7:0] layer0_N112_wire = {M0[121], M0[120], M0[95], M0[94], M0[59], M0[58], M0[47], M0[46]};
layer0_N112 layer0_N112_inst (.M0(layer0_N112_wire), .M1(M1[225:224]));

wire [7:0] layer0_N113_wire = {M0[113], M0[112], M0[81], M0[80], M0[79], M0[78], M0[49], M0[48]};
layer0_N113 layer0_N113_inst (.M0(layer0_N113_wire), .M1(M1[227:226]));

wire [7:0] layer0_N114_wire = {M0[69], M0[68], M0[51], M0[50], M0[35], M0[34], M0[1], M0[0]};
layer0_N114 layer0_N114_inst (.M0(layer0_N114_wire), .M1(M1[229:228]));

wire [7:0] layer0_N115_wire = {M0[113], M0[112], M0[83], M0[82], M0[71], M0[70], M0[61], M0[60]};
layer0_N115 layer0_N115_inst (.M0(layer0_N115_wire), .M1(M1[231:230]));

wire [7:0] layer0_N116_wire = {M0[113], M0[112], M0[61], M0[60], M0[57], M0[56], M0[41], M0[40]};
layer0_N116 layer0_N116_inst (.M0(layer0_N116_wire), .M1(M1[233:232]));

wire [7:0] layer0_N117_wire = {M0[123], M0[122], M0[59], M0[58], M0[53], M0[52], M0[33], M0[32]};
layer0_N117 layer0_N117_inst (.M0(layer0_N117_wire), .M1(M1[235:234]));

wire [7:0] layer0_N118_wire = {M0[81], M0[80], M0[59], M0[58], M0[49], M0[48], M0[21], M0[20]};
layer0_N118 layer0_N118_inst (.M0(layer0_N118_wire), .M1(M1[237:236]));

wire [7:0] layer0_N119_wire = {M0[91], M0[90], M0[85], M0[84], M0[57], M0[56], M0[13], M0[12]};
layer0_N119 layer0_N119_inst (.M0(layer0_N119_wire), .M1(M1[239:238]));

wire [7:0] layer0_N120_wire = {M0[99], M0[98], M0[69], M0[68], M0[65], M0[64], M0[13], M0[12]};
layer0_N120 layer0_N120_inst (.M0(layer0_N120_wire), .M1(M1[241:240]));

wire [7:0] layer0_N121_wire = {M0[123], M0[122], M0[103], M0[102], M0[65], M0[64], M0[35], M0[34]};
layer0_N121 layer0_N121_inst (.M0(layer0_N121_wire), .M1(M1[243:242]));

wire [7:0] layer0_N122_wire = {M0[69], M0[68], M0[65], M0[64], M0[17], M0[16], M0[3], M0[2]};
layer0_N122 layer0_N122_inst (.M0(layer0_N122_wire), .M1(M1[245:244]));

wire [7:0] layer0_N123_wire = {M0[105], M0[104], M0[97], M0[96], M0[59], M0[58], M0[23], M0[22]};
layer0_N123 layer0_N123_inst (.M0(layer0_N123_wire), .M1(M1[247:246]));

wire [7:0] layer0_N124_wire = {M0[113], M0[112], M0[95], M0[94], M0[67], M0[66], M0[47], M0[46]};
layer0_N124 layer0_N124_inst (.M0(layer0_N124_wire), .M1(M1[249:248]));

wire [7:0] layer0_N125_wire = {M0[81], M0[80], M0[57], M0[56], M0[29], M0[28], M0[13], M0[12]};
layer0_N125 layer0_N125_inst (.M0(layer0_N125_wire), .M1(M1[251:250]));

wire [7:0] layer0_N126_wire = {M0[95], M0[94], M0[31], M0[30], M0[21], M0[20], M0[3], M0[2]};
layer0_N126 layer0_N126_inst (.M0(layer0_N126_wire), .M1(M1[253:252]));

wire [7:0] layer0_N127_wire = {M0[123], M0[122], M0[79], M0[78], M0[69], M0[68], M0[31], M0[30]};
layer0_N127 layer0_N127_inst (.M0(layer0_N127_wire), .M1(M1[255:254]));

endmodule